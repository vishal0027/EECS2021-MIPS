module Engine(z, a, b);

output z;
input[1:0] a, b;

...

endmodule
 module rm(out, in1, in2);
  output out;
  input[1:0] in1, in2;
